`include "alu_intf.sv"
`include "alu_tx.sv"
`include "alu_gen.sv"
`include "alu_drv.sv"
`include "alu_mon.sv"
`include "alu_scb.sv"
`include "alu_cov.sv"
`include "alu_cfg.sv"
`include "alu_env.sv"
`include "alu_tb.sv"
`include "alu_top.sv"